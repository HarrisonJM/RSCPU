--OPLUT
-- Code your testbench here
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity OPLUT is
port( 
		addr: in std_logic_vector(6 downto 0);
		micCode_out: out std_logic_vector(18 downto 0)
    );
end entity;

architecture struct of OPLUT is

	type micMem is array (0 to 127) of std_logic_vector(18 downto 0);
	
	--0000 = uncondtional
	--0001 = Jump on Zero
	--0010 = Jump on !zero
	
	--0011 = Overflow 
	--0100 = !overflow
	
	--0101 = Carry
	--0110 = !Carry
	
	--0111 = Negative
	--1000 = !negative
	
	
	constant micCode : micMem := 
	( --GO THROUGH TABLE AND DOUBLE CHECK ALLL ENTRIES!!!
		--Cond	      BT 	 MicopAddr	NextAddress
	  0  => "0000" & "00" & "000000" & "0000001",     -- NOP
	  1  => "0000" & "00" & "000001" & "0000010",     -- FETCH1
	  2  => "0000" & "00" & "000010" & "0000011",     -- FETCH2
	  3  => "0000" & "01" & "000011" & "0000000",     -- FETCH3
	  
	  4  => "0000" & "10" & "000000" & "0111101",     -- LDAC0
	  5  => "0000" & "00" & "000100" & "0100001",     -- LDAC4
	  	  
	  8  => "0000" & "10" & "000000" & "0111101",     -- STAC0
	  9  => "0000" & "00" & "000101" & "0100010",     -- STAC4
	  
	  12 => "0000" & "00" & "000110" & "0000001",     -- MVAC1 
	  
	  16 => "0000" & "00" & "000111" & "0000001",     -- MOVR1
	  
	  20 => "0000" & "00" & "001000" & "0010101",     -- JUMP1
	  21 => "0000" & "00" & "001001" & "0010110",     -- JUMP2
	  22 => "0000" & "00" & "001010" & "0000001",     -- JUMP3

	  ----------------------------	  ----------------------------	  ----------------------------
	  24 => "0001" & "00" & "000000" & "0011001",     -- JMPZ1  --Jump if zero
	  25 => "0000" & "00" & "010001" & "0011010",     -- JMPZN1 --fail state
	  ---------------------------- 	 ----------------------------	  ----------------------------

	  26 => "0000" & "00" & "010001" & "0000001",     -- JMPF2 --Universal second fail state

	  28 => "0010" & "00" & "000000" & "0010100",     -- JPNZ1	 --Jump if not zero
 	  29 => "0000" & "00" & "010001" & "0011010",     -- JPNZN1 --fail state	 

	  32 => "0000" & "00" & "001101" & "0000001",     -- ADD1
	  33 => "0000" & "00" & "001011" & "0000001",     -- LDAC5
	  34 => "0000" & "00" & "001100" & "0000001",     -- STAC5

	  36 => "0000" & "00" & "001110" & "0000001",     -- SUB1
	  
	  40 => "0000" & "00" & "001111" & "0000001",     -- INAC1
	  
	  44 => "0000" & "00" & "010000" & "0000001",     -- CLAC1	  
	   
	  48 => "0000" & "00" & "010010" & "0000001",     -- AND1  
	  52 => "0000" & "00" & "010011" & "0000001",     -- OR1  
	  56 => "0000" & "00" & "010100" & "0000001",     -- XOR1  
	  60 => "0000" & "00" & "010101" & "0000001",     -- NOT1
	  	  
	  61 => "0000" & "00" & "010110" & "0111110",     -- SLSUB0
	  62 => "0000" & "00" & "010111" & "0111111",     -- SLSUB1
	  63 => "0000" & "11" & "011000" & "0000000",     -- SLSUB2
	  
	  64 => "0000" & "00" & "011110" & "1000001",     -- LDIND1
	  65 => "0000" & "00" & "000100" & "1000010",     -- LDIND2
	  66 => "0000" & "00" & "001011" & "0000001",     -- LDIND3
	  
	  68 => "0000" & "00" & "011110" & "1000101",     --STIND1	  
	  69 => "0000" & "00" & "000101" & "1000110",     --STIND2
	  70 => "0000" & "00" & "001100" & "0000001",     --STIND3
	  
	  72 => "0000" & "00" & "000101" & "1001001",     --LDINDAC1
	  73 => "0000" & "00" & "011111" & "1001010",     --LDINDAC2
	  74 => "0000" & "00" & "000101" & "1001011",     --LDINDAC3
	  75 => "0000" & "00" & "100000" & "0000001",     --LDINDAC4
	  
	  76 => "0000" & "00" & "011100" & "0000001",     -- INDD, decrement
	  
	  80 => "0000" & "00" & "011011" & "0000001",     -- INDIN
	  
	  84 => "0101" & "00" & "000000" & "0010100",     -- JMPC, jump on carry
	  85 => "0000" & "00" & "010001" & "0011010",     --Fail state
	  
	  88 => "0110" & "00" & "000000" & "0010100",     --JMPNC, jump on no carry
	  89 => "0000" & "00" & "010001" & "0011010",     --Fail state 
	  
	  92 => "0011" & "00" & "000000" & "0010100",     --JMPO Jump on OVerFlow
	  93 => "0000" & "00" & "010001" & "0011010",     --Fail state
	  
	  96 => "0100" & "00" & "000000" & "0010100",     --JPNO Jump on No Overflow
	  97 => "0000" & "00" & "010001" & "0011010",     --Fail state
	  
	  100 => "0111" & "00" & "000000" & "0010100",    --JMPN Jump on Negative
	  101 => "0000" & "00" & "010001" & "0011010",    --JMPNN Fail state
	  
	  104 => "1000" & "00" & "000000" & "0010100",    --JPNN Jump on No Negative
	  105 => "0000" & "00" & "010001" & "0011010",    --JPNNN Fail state
	  
	  108 => "0000" & "00" & "011101" & "0000001",    -- ADDC
	  
	  112 => "0000" & "00" & "011010" & "0000001",    --MVTI
 	  
 	  116 => "0000" & "00" & "011001" & "0000001",    --MVIT
	  
	  others => (others => '0')
	);

begin

	micCode_out <= micCode(to_integer(unsigned(addr)));


end struct;